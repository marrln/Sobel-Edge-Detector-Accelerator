library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use WORK.MY_TYPES.ALL;

entity manhattan_norm is
    port (
        clk     : in  std_logic;
        rst_n   : in  std_logic;
        s_valid : in  std_logic;
        s_ready : out std_logic;
        s_last  : in  std_logic;
        s_data  : in  gradient_pair;
        m_valid : out std_logic;
        m_ready : in  std_logic;
        m_last  : out std_logic;
        m_data  : out std_logic_vector(pixel_width - 1 downto 0)
    );
end entity manhattan_norm;

architecture Behavioral of manhattan_norm is
    signal abs_gx   : unsigned(gradient_width - 1 downto 0);
    signal abs_gy   : unsigned(gradient_width - 1 downto 0);
    signal sum_temp : unsigned(gradient_width downto 0);  -- one extra bit for carry
begin
    -- AXI handshake passthrough
    s_ready <= m_ready;
    m_valid <= s_valid;
    m_last  <= s_last;

    process(clk, rst_n)
    begin
        if rst_n = '0' then
            m_data   <= (others => '0');
            abs_gx   <= (others => '0');
            abs_gy   <= (others => '0');
            sum_temp <= (others => '0');

        elsif rising_edge(clk) then
            if m_ready = '1' then
                -- Compute absolute values using abs()
                abs_gx <= unsigned(abs(signed(s_data(0))));
                abs_gy <= unsigned(abs(signed(s_data(1))));

                -- Sum with one extra bit for carry
                sum_temp <= resize(abs_gx, sum_temp'length) + resize(abs_gy, sum_temp'length);

                -- Saturate to 8-bit pixel output
                if sum_temp > to_unsigned(255, sum_temp'length) then
                    m_data <= std_logic_vector(to_unsigned(255, pixel_width));
                else
                    m_data <= std_logic_vector(resize(sum_temp, pixel_width));
                end if;
            end if;
        end if;
    end process;
end Behavioral;
